library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity project_tb is
end project_tb;

architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 100 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst	                : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		        : std_logic := '0';
signal   mem_o_data,mem_i_data	: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		        : std_logic;
signal   update_addr            : std_logic_vector(15 downto 0);
signal   update_mem             : std_logic;
signal   new_ind               : std_logic_vector(7 downto 0);

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);

-- come da esempio su specifica
signal RAM: ram_type := (0 => std_logic_vector(to_unsigned( 7 , 8)),
                         1 => std_logic_vector(to_unsigned( 23 , 8)),
                         2 => std_logic_vector(to_unsigned( 80 , 8)),
                         3 => std_logic_vector(to_unsigned( 29 , 8)),
                         4 => std_logic_vector(to_unsigned( 1 , 8)),
                         5 => std_logic_vector(to_unsigned( 57 , 8)),
                         6 => std_logic_vector(to_unsigned( 48 , 8)),
                         7 => std_logic_vector(to_unsigned( 112 , 8)),
                         8 => std_logic_vector(to_unsigned( 48 , 8)),
			 others => (others =>'0'));

component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_start       : in  std_logic;
      i_rst         : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            elsif update_mem = '1' then
                RAM(conv_integer(update_addr)) <= new_ind;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end process;


test : process is
begin
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    tb_start <= '1';
    wait for 1000 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    update_addr <= "0000000000001000";
    new_ind <= std_logic_vector(to_unsigned(49, 8));
    update_mem <= '1';
    wait for 200 ns;

    if RAM(9) = std_logic_vector(to_unsigned(  225, 8)) then
        report "PRIMO TEST PASSATO";
    else
        report "PRIMO TEST FALLITO, found " & integer'image(to_integer(unsigned(RAM(9))));
    end if;
    wait for c_CLOCK_PERIOD;
    update_mem <= '0';
    tb_start <= '1';
    report "MEM aggiornata " & integer'image(to_integer(unsigned(RAM(8))));
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    
    wait for 100 ns;
    update_addr <= "0000000000001000";
        new_ind <= std_logic_vector(to_unsigned(50, 8));
        update_mem <= '1';
        wait for 200 ns;
    
        if RAM(9) = std_logic_vector(to_unsigned(  226, 8)) then
            report "SECONDO TEST PASSATO";
        else
            report "SECONDO TEST FALLITO, found " & integer'image(to_integer(unsigned(RAM(9))));
        end if;
        wait for c_CLOCK_PERIOD;
        update_mem <= '0';
        tb_start <= '1';
        report "MEM aggiornata " & integer'image(to_integer(unsigned(RAM(8))));
        wait for c_CLOCK_PERIOD;
        wait until tb_done = '1';
        wait for c_CLOCK_PERIOD;
        tb_start <= '0';
        wait until tb_done = '0';
        
         wait for 100 ns;
           update_addr <= "0000000000001000";
               new_ind <= std_logic_vector(to_unsigned(51, 8));
               update_mem <= '1';
               wait for 200 ns;
           
               if RAM(9) = std_logic_vector(to_unsigned(  228, 8)) then
                   report "TERZO TEST PASSATO";
               else
                   report "TERZO TEST FALLITO, found " & integer'image(to_integer(unsigned(RAM(9))));
               end if;
               wait for c_CLOCK_PERIOD;
               update_mem <= '0';
               
               --blocco di reset 
               wait for 100 ns;
                   wait for c_CLOCK_PERIOD;
                   tb_rst <= '1';
                   wait for c_CLOCK_PERIOD;
                   tb_rst <= '0';
                   wait for c_CLOCK_PERIOD;
                   tb_start <= '1';
                   wait for 1000 ns;
                   wait for c_CLOCK_PERIOD;
                   tb_rst <= '1';
                   wait for c_CLOCK_PERIOD;
                   tb_rst <= '0';
                   wait for 200 ns; 
                   wait for c_CLOCK_PERIOD;
                                      tb_rst <= '1';
                                      wait for c_CLOCK_PERIOD;
                                      tb_rst <= '0';
                                      wait for c_CLOCK_PERIOD;
                                      tb_start <= '1';
                                      wait for 1000 ns;
                                      wait for c_CLOCK_PERIOD;
                                      tb_rst <= '1';
                                      wait for c_CLOCK_PERIOD;
                                      tb_rst <= '0';
                                      wait for 200 ns; 
                                      wait for c_CLOCK_PERIOD;
                                                         tb_rst <= '1';
                                                         wait for c_CLOCK_PERIOD;
                                                         tb_rst <= '0';
                                                         wait for c_CLOCK_PERIOD;
                                                         tb_start <= '1';
                                                         wait for 1000 ns;
                                                         wait for c_CLOCK_PERIOD;
                                                         tb_rst <= '1';
                                                         wait for c_CLOCK_PERIOD;
                                                         tb_rst <= '0';
                                                         wait for 200 ns; 
                   
                   
               tb_start <= '1';
               report "MEM aggiornata " & integer'image(to_integer(unsigned(RAM(8))));
               wait for c_CLOCK_PERIOD;
               wait until tb_done = '1';
               wait for c_CLOCK_PERIOD;
               tb_start <= '0';
               wait until tb_done = '0';
    
                        wait for 100 ns;
                          update_addr <= "0000000000001000";
                              new_ind <= std_logic_vector(to_unsigned(52, 8));
                              update_mem <= '1';
                              wait for 200 ns;
                          
                              if RAM(9) = std_logic_vector(to_unsigned(  232, 8)) then
                                  report "QUARTO TEST PASSATO";
                              else
                                  report "QUARTO TEST FALLITO, found " & integer'image(to_integer(unsigned(RAM(9))));
                              end if;
                              wait for c_CLOCK_PERIOD;
                              update_mem <= '0';
                              tb_start <= '1';
                              report "MEM aggiornata " & integer'image(to_integer(unsigned(RAM(8))));
                              wait for c_CLOCK_PERIOD;
                              wait until tb_done = '1';
                              wait for c_CLOCK_PERIOD;
                              tb_start <= '0';
                              wait until tb_done = '0';
    wait for 100 ns;
    

    -- Maschera di output = 1 - 110 - 1000
    assert RAM(9) = std_logic_vector(to_unsigned( 52 , 8)) report "QUINTO TEST FALLITO. Expected  130  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

    assert false report "Simulation Ended!, QUINTO TEST PASSATO" severity failure;
end process test;

end projecttb; 
